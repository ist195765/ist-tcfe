.OP
Vs 1 0 0.0 AC 1.0 sin(0 1 1000)
R1 1 2 1.013609e+03 
R2 3 2 2.016578e+03 
R3 2 5 3.006816e+03 
R4 5 0 4.049229e+03 
R5 5 6 3.053925e+03 
R6 9 7 2.092502e+03 
R7 7 8 1.022320e+03 
C1 6 8 1.029587e-06 
.IC v(6) = 5.853598e+00 v(8) = -2.978754e+00
Vaux 0 9 0.000000e+00 
Hd 5 8 Vaux 8.321035e+03 
Gb 6 3 (2,5) 7.213324e-03 
.END
